VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO non_hwt
  CLASS BLOCK ;
  FOREIGN non_hwt ;
  ORIGIN 3.500 -0.400 ;
  SIZE 31.000 BY 21.200 ;
  PIN A
    PORT
      LAYER metal1 ;
        RECT 4.400 7.600 5.200 10.400 ;
      LAYER metal2 ;
        RECT 4.400 7.600 5.200 8.400 ;
        RECT 4.500 6.400 5.100 7.600 ;
        RECT 4.400 5.600 5.200 6.400 ;
      LAYER metal3 ;
        RECT 4.400 6.300 5.200 6.400 ;
        RECT -3.500 5.700 5.200 6.300 ;
        RECT 4.400 5.600 5.200 5.700 ;
    END
  END A
  PIN B
    PORT
      LAYER metal1 ;
        RECT -2.000 14.300 -1.200 14.400 ;
        RECT 1.200 14.300 2.000 15.200 ;
        RECT -2.000 13.700 2.000 14.300 ;
        RECT -2.000 13.600 -1.200 13.700 ;
        RECT 1.200 13.600 2.000 13.700 ;
      LAYER metal2 ;
        RECT -2.000 13.600 -1.200 14.400 ;
      LAYER metal3 ;
        RECT -2.000 14.300 -1.200 14.400 ;
        RECT -3.500 13.700 -1.200 14.300 ;
        RECT -2.000 13.600 -1.200 13.700 ;
    END
  END B
  PIN C
    PORT
      LAYER metal1 ;
        RECT 18.800 15.600 19.600 17.200 ;
      LAYER metal2 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 18.900 10.400 19.500 15.600 ;
        RECT 18.800 9.600 19.600 10.400 ;
      LAYER metal3 ;
        RECT 18.800 10.300 19.600 10.400 ;
        RECT 18.800 9.700 27.500 10.300 ;
        RECT 18.800 9.600 19.600 9.700 ;
    END
  END C
  PIN D
    PORT
      LAYER metal1 ;
        RECT 22.000 16.300 22.800 17.200 ;
        RECT 23.600 16.300 24.400 16.400 ;
        RECT 22.000 15.700 24.400 16.300 ;
        RECT 22.000 15.600 22.800 15.700 ;
        RECT 23.600 15.600 24.400 15.700 ;
      LAYER metal2 ;
        RECT 23.600 15.600 24.400 16.400 ;
        RECT 23.700 6.400 24.300 15.600 ;
        RECT 23.600 5.600 24.400 6.400 ;
      LAYER metal3 ;
        RECT 23.600 6.300 24.400 6.400 ;
        RECT 23.600 5.700 27.500 6.300 ;
        RECT 23.600 5.600 24.400 5.700 ;
    END
  END D
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 6.000 12.400 6.800 19.800 ;
        RECT 6.000 10.200 6.600 12.400 ;
        RECT 6.000 2.200 6.800 10.200 ;
      LAYER via1 ;
        RECT 6.000 13.600 6.800 14.400 ;
      LAYER metal2 ;
        RECT 6.000 13.600 6.800 14.400 ;
        RECT 6.100 10.400 6.700 13.600 ;
        RECT 6.000 9.600 6.800 10.400 ;
      LAYER metal3 ;
        RECT 6.000 10.300 6.800 10.400 ;
        RECT -3.500 9.700 6.800 10.300 ;
        RECT 6.000 9.600 6.800 9.700 ;
    END
  END Y
  OBS
      LAYER metal1 ;
        RECT 0.400 20.400 23.600 21.600 ;
        RECT 1.200 15.800 2.000 20.400 ;
        RECT 3.800 16.400 4.600 19.800 ;
        RECT 2.800 15.800 4.600 16.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 2.800 12.300 3.600 15.800 ;
        RECT 9.200 15.200 10.000 19.800 ;
        RECT 11.400 15.800 12.200 20.400 ;
        RECT 14.000 15.800 14.800 19.800 ;
        RECT 15.600 17.800 16.400 20.400 ;
        RECT 15.400 16.400 16.200 17.200 ;
        RECT 7.800 14.600 10.000 15.200 ;
        RECT 4.400 12.300 5.200 12.400 ;
        RECT 2.800 11.700 5.200 12.300 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 2.800 2.200 3.600 11.700 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 7.800 11.600 8.400 14.600 ;
        RECT 9.200 11.600 10.000 13.200 ;
        RECT 12.400 12.800 13.200 14.400 ;
        RECT 14.000 12.400 14.600 15.800 ;
        RECT 15.600 15.600 16.400 16.400 ;
        RECT 15.600 14.300 16.400 14.400 ;
        RECT 17.200 14.300 18.000 19.800 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 15.600 13.700 18.000 14.300 ;
        RECT 15.600 13.600 16.400 13.700 ;
        RECT 10.800 12.200 11.600 12.400 ;
        RECT 14.000 12.200 14.800 12.400 ;
        RECT 15.600 12.200 16.400 12.400 ;
        RECT 10.800 11.600 12.400 12.200 ;
        RECT 14.000 11.600 16.400 12.200 ;
        RECT 7.200 10.800 8.400 11.600 ;
        RECT 11.600 11.200 12.400 11.600 ;
        RECT 7.800 10.200 8.400 10.800 ;
        RECT 15.600 10.200 16.200 11.600 ;
        RECT 7.800 9.600 10.000 10.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 9.000 ;
        RECT 9.200 2.200 10.000 9.600 ;
        RECT 10.800 9.600 14.800 10.200 ;
        RECT 10.800 2.200 11.600 9.600 ;
        RECT 12.400 1.600 13.200 9.000 ;
        RECT 14.000 2.200 14.800 9.600 ;
        RECT 15.600 2.200 16.400 10.200 ;
        RECT 17.200 2.200 18.000 13.700 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 20.400 2.200 21.200 19.800 ;
        RECT 22.000 17.800 22.800 20.400 ;
        RECT 22.000 1.600 22.800 6.200 ;
        RECT 0.400 0.400 23.600 1.600 ;
      LAYER via1 ;
        RECT 12.400 13.600 13.200 14.400 ;
        RECT 20.400 15.600 21.200 16.400 ;
      LAYER metal2 ;
        RECT 15.600 15.600 16.400 16.400 ;
        RECT 20.400 15.600 21.200 16.400 ;
        RECT 12.400 13.600 13.200 14.400 ;
        RECT 15.600 13.600 16.400 14.400 ;
        RECT 4.400 11.600 5.200 12.400 ;
        RECT 9.200 11.600 10.000 12.400 ;
        RECT 10.800 11.600 11.600 12.400 ;
        RECT 14.000 11.600 14.800 12.400 ;
        RECT 9.300 10.400 9.900 11.600 ;
        RECT 14.100 10.400 14.700 11.600 ;
        RECT 9.200 9.600 10.000 10.400 ;
        RECT 14.000 9.600 14.800 10.400 ;
      LAYER metal3 ;
        RECT 15.600 16.300 16.400 16.400 ;
        RECT 20.400 16.300 21.200 16.400 ;
        RECT 15.600 15.700 21.200 16.300 ;
        RECT 15.600 15.600 16.400 15.700 ;
        RECT 20.400 15.600 21.200 15.700 ;
        RECT 12.400 14.300 13.200 14.400 ;
        RECT 15.600 14.300 16.400 14.400 ;
        RECT 12.400 13.700 16.400 14.300 ;
        RECT 12.400 13.600 13.200 13.700 ;
        RECT 15.600 13.600 16.400 13.700 ;
        RECT 4.400 12.300 5.200 12.400 ;
        RECT 10.800 12.300 11.600 12.400 ;
        RECT 4.400 11.700 11.600 12.300 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 10.800 11.600 11.600 11.700 ;
        RECT 9.200 10.300 10.000 10.400 ;
        RECT 14.000 10.300 14.800 10.400 ;
        RECT 9.200 9.700 14.800 10.300 ;
        RECT 9.200 9.600 10.000 9.700 ;
        RECT 14.000 9.600 14.800 9.700 ;
  END
END non_hwt
END LIBRARY


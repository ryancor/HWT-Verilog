VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hwt
  CLASS BLOCK ;
  FOREIGN hwt ;
  ORIGIN 3.500 1.000 ;
  SIZE 51.800 BY 27.300 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 20.400 44.400 21.600 ;
        RECT 1.200 15.800 2.000 20.400 ;
        RECT 6.000 13.800 6.800 20.400 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 22.600 15.800 23.400 20.400 ;
        RECT 26.800 17.800 27.600 20.400 ;
        RECT 38.000 15.800 38.800 20.400 ;
        RECT 41.200 15.800 42.000 20.400 ;
      LAYER via1 ;
        RECT 27.500 20.600 28.300 21.400 ;
        RECT 28.500 20.600 29.300 21.400 ;
        RECT 29.500 20.600 30.300 21.400 ;
        RECT 30.500 20.600 31.300 21.400 ;
        RECT 31.500 20.600 32.300 21.400 ;
        RECT 32.500 20.600 33.300 21.400 ;
      LAYER metal2 ;
        RECT 29.800 21.400 31.000 21.600 ;
        RECT 27.500 20.600 33.300 21.400 ;
        RECT 29.800 20.400 31.000 20.600 ;
      LAYER via2 ;
        RECT 28.500 20.600 29.300 21.400 ;
        RECT 29.500 20.600 30.300 21.400 ;
        RECT 30.500 20.600 31.300 21.400 ;
        RECT 31.500 20.600 32.300 21.400 ;
        RECT 32.500 20.600 33.300 21.400 ;
      LAYER metal3 ;
        RECT 27.400 20.400 33.400 21.600 ;
      LAYER via3 ;
        RECT 27.600 20.600 28.400 21.400 ;
        RECT 28.800 20.600 29.600 21.400 ;
        RECT 30.000 20.600 30.800 21.400 ;
        RECT 31.200 20.600 32.000 21.400 ;
        RECT 32.400 20.600 33.200 21.400 ;
      LAYER metal4 ;
        RECT 27.200 -1.000 33.600 21.600 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 6.000 1.600 6.800 6.200 ;
        RECT 9.200 1.600 10.000 5.800 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 23.600 1.600 24.400 9.000 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 38.000 1.600 38.800 6.200 ;
        RECT 41.200 1.600 42.000 9.000 ;
        RECT 0.400 0.400 44.400 1.600 ;
      LAYER via1 ;
        RECT 11.500 0.600 12.300 1.400 ;
        RECT 12.500 0.600 13.300 1.400 ;
        RECT 13.500 0.600 14.300 1.400 ;
        RECT 14.500 0.600 15.300 1.400 ;
        RECT 15.500 0.600 16.300 1.400 ;
        RECT 16.500 0.600 17.300 1.400 ;
      LAYER metal2 ;
        RECT 13.800 1.400 15.000 1.600 ;
        RECT 11.500 0.600 17.300 1.400 ;
        RECT 13.800 0.400 15.000 0.600 ;
      LAYER via2 ;
        RECT 12.500 0.600 13.300 1.400 ;
        RECT 13.500 0.600 14.300 1.400 ;
        RECT 14.500 0.600 15.300 1.400 ;
        RECT 15.500 0.600 16.300 1.400 ;
        RECT 16.500 0.600 17.300 1.400 ;
      LAYER metal3 ;
        RECT 11.400 0.400 17.400 1.600 ;
      LAYER via3 ;
        RECT 11.600 0.600 12.400 1.400 ;
        RECT 12.800 0.600 13.600 1.400 ;
        RECT 14.000 0.600 14.800 1.400 ;
        RECT 15.200 0.600 16.000 1.400 ;
        RECT 16.400 0.600 17.200 1.400 ;
      LAYER metal4 ;
        RECT 11.200 -1.000 17.600 21.600 ;
    END
  END vdd
  PIN A
    PORT
      LAYER metal1 ;
        RECT 7.600 11.600 9.200 12.400 ;
        RECT 4.400 8.300 5.200 10.400 ;
        RECT 7.600 8.300 8.400 8.400 ;
        RECT 4.400 7.700 8.400 8.300 ;
        RECT 7.600 7.600 8.400 7.700 ;
      LAYER metal2 ;
        RECT 7.600 11.600 8.400 12.400 ;
        RECT 7.700 8.400 8.300 11.600 ;
        RECT 7.600 7.600 8.400 8.400 ;
        RECT 7.700 6.400 8.300 7.600 ;
        RECT 7.600 5.600 8.400 6.400 ;
      LAYER metal3 ;
        RECT 7.600 6.300 8.400 6.400 ;
        RECT -3.500 5.700 8.400 6.300 ;
        RECT 7.600 5.600 8.400 5.700 ;
    END
  END A
  PIN B
    PORT
      LAYER metal1 ;
        RECT 1.200 13.600 2.000 15.200 ;
        RECT 6.000 9.600 6.800 11.200 ;
      LAYER metal2 ;
        RECT 1.200 13.600 2.000 14.400 ;
        RECT 1.300 10.400 1.900 13.600 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 6.000 9.600 6.800 10.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT 6.000 10.300 6.800 10.400 ;
        RECT -3.500 9.700 6.800 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
        RECT 6.000 9.600 6.800 9.700 ;
    END
  END B
  PIN C
    PORT
      LAYER metal1 ;
        RECT 18.800 15.600 19.600 17.200 ;
        RECT 9.200 7.600 10.000 9.200 ;
      LAYER metal2 ;
        RECT 18.900 25.700 21.100 26.300 ;
        RECT 18.900 16.400 19.500 25.700 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 18.900 12.400 19.500 15.600 ;
        RECT 9.200 11.600 10.000 12.400 ;
        RECT 18.800 11.600 19.600 12.400 ;
        RECT 9.300 8.400 9.900 11.600 ;
        RECT 9.200 7.600 10.000 8.400 ;
      LAYER metal3 ;
        RECT 9.200 12.300 10.000 12.400 ;
        RECT 18.800 12.300 19.600 12.400 ;
        RECT 9.200 11.700 19.600 12.300 ;
        RECT 9.200 11.600 10.000 11.700 ;
        RECT 18.800 11.600 19.600 11.700 ;
    END
  END C
  PIN D
    PORT
      LAYER metal1 ;
        RECT 38.000 13.600 38.800 15.200 ;
      LAYER metal2 ;
        RECT 38.000 14.300 38.800 14.400 ;
        RECT 38.000 13.700 40.300 14.300 ;
        RECT 38.000 13.600 38.800 13.700 ;
        RECT 39.700 10.400 40.300 13.700 ;
        RECT 39.600 9.600 40.400 10.400 ;
      LAYER metal3 ;
        RECT 39.600 10.300 40.400 10.400 ;
        RECT 39.600 9.700 48.300 10.300 ;
        RECT 39.600 9.600 40.400 9.700 ;
    END
  END D
  PIN Y
    PORT
      LAYER metal1 ;
        RECT 42.800 12.400 43.600 19.800 ;
        RECT 43.000 10.200 43.600 12.400 ;
        RECT 42.800 6.300 43.600 10.200 ;
        RECT 44.400 6.300 45.200 6.400 ;
        RECT 42.800 5.700 45.200 6.300 ;
        RECT 42.800 2.200 43.600 5.700 ;
        RECT 44.400 5.600 45.200 5.700 ;
      LAYER metal2 ;
        RECT 44.400 5.600 45.200 6.400 ;
      LAYER metal3 ;
        RECT 44.400 6.300 45.200 6.400 ;
        RECT 44.400 5.700 48.300 6.300 ;
        RECT 44.400 5.600 45.200 5.700 ;
    END
  END Y
  OBS
      LAYER metal1 ;
        RECT 3.800 16.400 4.600 19.800 ;
        RECT 2.800 15.800 4.600 16.400 ;
        RECT 2.800 14.300 3.600 15.800 ;
        RECT 4.400 14.300 5.200 14.400 ;
        RECT 2.800 13.700 5.200 14.300 ;
        RECT 9.600 14.200 10.400 19.800 ;
        RECT 9.600 13.800 11.400 14.200 ;
        RECT 2.800 2.200 3.600 13.700 ;
        RECT 4.400 13.600 5.200 13.700 ;
        RECT 9.800 13.600 11.400 13.800 ;
        RECT 10.800 10.400 11.400 13.600 ;
        RECT 20.400 12.300 21.200 19.800 ;
        RECT 25.200 15.800 26.000 19.800 ;
        RECT 26.600 16.400 27.400 17.200 ;
        RECT 35.400 16.400 36.200 19.800 ;
        RECT 26.800 16.300 27.600 16.400 ;
        RECT 35.400 16.300 37.200 16.400 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 23.600 14.300 24.400 14.400 ;
        RECT 22.000 13.700 24.400 14.300 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 23.600 12.800 24.400 13.700 ;
        RECT 22.000 12.300 22.800 12.400 ;
        RECT 20.400 12.200 22.800 12.300 ;
        RECT 25.200 12.200 25.800 15.800 ;
        RECT 26.800 15.700 37.200 16.300 ;
        RECT 26.800 15.600 27.600 15.700 ;
        RECT 26.800 12.200 27.600 12.400 ;
        RECT 20.400 11.700 23.600 12.200 ;
        RECT 10.800 10.300 11.600 10.400 ;
        RECT 18.800 10.300 19.600 10.400 ;
        RECT 10.800 9.700 19.600 10.300 ;
        RECT 10.800 9.600 11.600 9.700 ;
        RECT 18.800 9.600 19.600 9.700 ;
        RECT 10.800 7.000 11.400 9.600 ;
        RECT 7.800 6.400 11.400 7.000 ;
        RECT 7.800 6.200 8.400 6.400 ;
        RECT 7.600 2.200 8.400 6.200 ;
        RECT 10.800 6.200 11.400 6.400 ;
        RECT 10.800 2.200 11.600 6.200 ;
        RECT 20.400 2.200 21.200 11.700 ;
        RECT 22.000 11.600 23.600 11.700 ;
        RECT 25.200 11.600 27.600 12.200 ;
        RECT 22.800 11.200 23.600 11.600 ;
        RECT 26.800 10.200 27.400 11.600 ;
        RECT 22.000 9.600 26.000 10.200 ;
        RECT 22.000 2.200 22.800 9.600 ;
        RECT 25.200 2.200 26.000 9.600 ;
        RECT 26.800 2.200 27.600 10.200 ;
        RECT 34.800 8.800 35.600 10.400 ;
        RECT 36.400 2.200 37.200 15.700 ;
        RECT 39.600 15.200 40.400 19.800 ;
        RECT 39.600 14.600 41.800 15.200 ;
        RECT 38.000 12.300 38.800 12.400 ;
        RECT 39.600 12.300 40.400 13.200 ;
        RECT 38.000 11.700 40.400 12.300 ;
        RECT 38.000 11.600 38.800 11.700 ;
        RECT 39.600 11.600 40.400 11.700 ;
        RECT 41.200 11.600 41.800 14.600 ;
        RECT 41.200 10.800 42.400 11.600 ;
        RECT 41.200 10.200 41.800 10.800 ;
        RECT 39.600 9.600 41.800 10.200 ;
        RECT 39.600 2.200 40.400 9.600 ;
      LAYER via1 ;
        RECT 26.800 11.600 27.600 12.400 ;
        RECT 34.800 9.600 35.600 10.400 ;
      LAYER metal2 ;
        RECT 4.400 13.600 5.200 14.400 ;
        RECT 22.000 13.600 22.800 14.400 ;
        RECT 26.800 11.600 27.600 12.400 ;
        RECT 38.000 11.600 38.800 12.400 ;
        RECT 18.800 9.600 19.600 10.400 ;
        RECT 34.800 9.600 35.600 10.400 ;
      LAYER metal3 ;
        RECT 4.400 14.300 5.200 14.400 ;
        RECT 22.000 14.300 22.800 14.400 ;
        RECT 4.400 13.700 22.800 14.300 ;
        RECT 4.400 13.600 5.200 13.700 ;
        RECT 22.000 13.600 22.800 13.700 ;
        RECT 26.800 12.300 27.600 12.400 ;
        RECT 38.000 12.300 38.800 12.400 ;
        RECT 26.800 11.700 38.800 12.300 ;
        RECT 26.800 11.600 27.600 11.700 ;
        RECT 38.000 11.600 38.800 11.700 ;
        RECT 18.800 10.300 19.600 10.400 ;
        RECT 34.800 10.300 35.600 10.400 ;
        RECT 18.800 9.700 35.600 10.300 ;
        RECT 18.800 9.600 19.600 9.700 ;
        RECT 34.800 9.600 35.600 9.700 ;
  END
END hwt
END LIBRARY

